----------------------------------------------------------------------------------
-- Engineer: Evan Votta
-- 
-- Design Name: 	Mips32 in VHDL
-- Module Name:   op_fetch - Behavioral 
-- Project Name: 	Mips32 in VHDL

-- Description: 	This file is used to simulate the data memory.
--
--						As you will notice, I like to capitalize keywords sometimes, a habit I
--						picked up from using SQL.
--
--						I'm used to documenting/commenting in a Javadoc style, I wasn't sure
--						if	there was a sort of standardized or common commenting style in VHDL. I saw
--						something like it in Verilog, but I figured if anything, the commenting
--						style would be more like Ada than C. From what I've read, Verilog is a bit
--						easier to learn, but it is for Software Developers pretending to be Logic
--						Design Engineers. VHDL is more exact, more precise, the engineer has better
--						command of what goes on in the design, so I guess I'm glad we learned VHDL
--						instead of Verilog. I hope you approve of the way I comment, I tried to make
--						it as descriptive as possible.
--
--						I also like to tab some lines out so that they are equal length and broken
--						down into sections, I picked up the habit writing assembly code for PIC16's.
--
----------------------------------------------------------------------------------
LIBRARY 	IEEE								;
	USE 	IEEE.STD_LOGIC_1164.ALL		;
	USE 	IEEE.STD_LOGIC_ARITH.ALL	;
	USE 	IEEE.STD_LOGIC_SIGNED.ALL	;



ENTITY data_memory IS
	PORT(
			-- First the inputs
			CLOCK 		: IN STD_LOGIC								;
			RESET 		: IN STD_LOGIC								;
			addr 			: IN STD_LOGIC_VECTOR (7 DOWNTO 0)	;
			write_data 	: IN STD_LOGIC_VECTOR (7 DOWNTO 0)	;
			mem_read 	: IN STD_LOGIC								;
			mem_write 	: IN STD_LOGIC								;
					
			-- Next the outputs (only one here)
			read_data 	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
		);
			
END data_memory;

ARCHITECTURE Behavioral OF data_memory IS

	-- Set the data slots, sizes, etc, etc.
   CONSTANT size 			: natural := 1024														;
   CONSTANT first_word 	: natural := 268500992												;
   CONSTANT last_word 	: natural := 268502015												;  
   TYPE 		mem_type IS ARRAY(natural range <>) OF std_logic_vector(31 DOWNTO 0)	;
   CONSTANT nod 			: std_logic_vector(31 downto 0) := (others => '0')			;
   
	
	
	-- Memory words --
   CONSTANT data_at_init : mem_type(0 to size-1) :=   
		(
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000010011",
			"00100000011101110110111101001000",	"01111001011011100110000101101101",
			"01100010011010010100011000100000",	"01100011011000010110111001101111",
			"01101110001000000110100101100011",	"01100101011000100110110101110101",
			"01110100001000000111001101110010",	"01100101011001110010000001101111",
			"01100001011100100110010101101110",	"00100000001111110110010101110100",
			"00111100001000000011001000101000",	"00100000011110000010000000111101",
			"00110001001000000011110100111100",	"00100000000000000010100100111001",
			"01100101011010000101010000000000",	"01100010011010010100011000100000",
			"01100011011000010110111001101111",	"01101110001000000110100101100011",
			"01100101011000100110110101110101",	"01100001001000000111001101110010",
			"00001010001110100110010101110010",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000", "00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000",
			"00000000000000000000000000000000",	"00000000000000000000000000000000"
	);
	-- end memory words, obviously --

   -- Internal signal declarations
   SIGNAL mem : mem_type(first_word TO last_word);
	
	BEGIN
		-- begin
	
		run : PROCESS (CLOCK, RESET)
			-- start process
			BEGIN
				-- Begin
			
				-- IF 1 --
				IF(RESET ='1') 							THEN
						mem(first_word 			TO first_word+size-1) 	<= data_at_init	;
						mem(first_word+size-1 	TO last_word		  ) 	<= (others=>nod)	;
				-- END IF 1 --
						
				-- IF 2 --
				ELSIF (CLOCK'EVENT AND CLOCK = '1') 
						AND (mem_write = '1') THEN
					mem(conv_integer(unsigned(addr))) 					<= write_data		;
				END IF;
				-- END IF @ --
	
	
		END PROCESS run;
		-- END the process : run --
		
	read_data <= mem(conv_integer(unsigned(addr)))
		WHEN (mem_read = '1')
		ELSE nod;

END Behavioral;